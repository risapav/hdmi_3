//App app(.pixel_clk(clk_25), .pixel_clk10(clk_250), .clk(clk_32));

module App (pixel_clk, pixel_clk10, clk);

input wire	pixel_clk, pixel_clk10, clk;



endmodule